
module FIFO_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] DIFF;
  input CI;
  output CO;
  wire   n3, n4, n6, n8, n9, n10, n11, n12, n13, n15, n17, n18, n19, n20, n21,
         n22, n23, n24, n47, n48, n49, n50;

  NAND2X1 U8 ( .A(A[1]), .B(n50), .Y(n10) );
  NOR2X1 U9 ( .A(A[1]), .B(n50), .Y(n11) );
  NAND2X1 U11 ( .A(n10), .B(n6), .Y(n21) );
  OAI21X1 U12 ( .A(n9), .B(n11), .C(n10), .Y(n12) );
  XOR2X1 U13 ( .A(n21), .B(n9), .Y(DIFF[1]) );
  NAND2X1 U14 ( .A(A[2]), .B(n3), .Y(n13) );
  NAND2X1 U17 ( .A(n13), .B(n48), .Y(n22) );
  AOI21X1 U20 ( .A(n48), .B(n12), .C(n15), .Y(n17) );
  XNOR2X1 U21 ( .A(n47), .B(n22), .Y(DIFF[2]) );
  NAND2X1 U22 ( .A(A[3]), .B(n4), .Y(n18) );
  NOR2X1 U23 ( .A(A[3]), .B(n4), .Y(n19) );
  NAND2X1 U25 ( .A(n18), .B(n8), .Y(n23) );
  OAI21X1 U26 ( .A(n19), .B(n17), .C(n18), .Y(n20) );
  XOR2X1 U27 ( .A(n17), .B(n23), .Y(DIFF[3]) );
  XOR2X1 U29 ( .A(n20), .B(n24), .Y(DIFF[4]) );
  INVX2 U33 ( .A(B[1]), .Y(n50) );
  OAI21X1 U34 ( .A(n9), .B(n11), .C(n10), .Y(n47) );
  XNOR2X1 U35 ( .A(B[4]), .B(A[4]), .Y(n24) );
  INVX2 U36 ( .A(A[0]), .Y(n49) );
  XOR2X1 U37 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
  OR2X2 U38 ( .A(A[2]), .B(n3), .Y(n48) );
  AND2X2 U39 ( .A(n49), .B(B[0]), .Y(n9) );
  INVX2 U40 ( .A(n19), .Y(n8) );
  INVX2 U41 ( .A(n11), .Y(n6) );
  INVX2 U42 ( .A(B[3]), .Y(n4) );
  INVX2 U43 ( .A(B[2]), .Y(n3) );
  INVX2 U44 ( .A(n13), .Y(n15) );
endmodule


module FIFO_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry_4_), .B(A[4]), .Y(SUM[4]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry_4_), .B(A[4]), .Y(SUM[4]) );
endmodule


module FIFO ( clk, reset, data_in, put, get, data_out, fillcount, empty, full
 );
  input [7:0] data_in;
  output [7:0] data_out;
  output [4:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   n11, n12, n13, n14, rd_ptr_4_, n33, n34, n35, n36, n37, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n365, n368, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n697, n698, n699, n700, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, SYNOPSYS_UNCONNECTED_1;
  wire   [4:0] wr_ptr;
  wire   [127:0] fifo;

  DFFPOSX1 rd_ptr_reg_0_ ( .D(n1057), .CLK(clk), .Q(n11) );
  DFFPOSX1 data_out_reg_7_ ( .D(n1058), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n1059), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n1060), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n1061), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n1062), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n1063), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n1064), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n1065), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n1066), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n1067), .CLK(clk), .Q(n12) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n1068), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n1069), .CLK(clk), .Q(rd_ptr_4_) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n700), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 wr_ptr_reg_0_ ( .D(n699), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n698), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n697), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n1070), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 fifo_reg_3__7_ ( .D(n695), .CLK(clk), .Q(fifo[31]) );
  DFFPOSX1 fifo_reg_3__5_ ( .D(n694), .CLK(clk), .Q(fifo[29]) );
  DFFPOSX1 fifo_reg_3__3_ ( .D(n693), .CLK(clk), .Q(fifo[27]) );
  DFFPOSX1 fifo_reg_3__1_ ( .D(n692), .CLK(clk), .Q(fifo[25]) );
  DFFPOSX1 fifo_reg_3__0_ ( .D(n691), .CLK(clk), .Q(fifo[24]) );
  DFFPOSX1 fifo_reg_3__2_ ( .D(n690), .CLK(clk), .Q(fifo[26]) );
  DFFPOSX1 fifo_reg_3__4_ ( .D(n689), .CLK(clk), .Q(fifo[28]) );
  DFFPOSX1 fifo_reg_3__6_ ( .D(n688), .CLK(clk), .Q(fifo[30]) );
  DFFPOSX1 fifo_reg_2__7_ ( .D(n687), .CLK(clk), .Q(fifo[23]) );
  DFFPOSX1 fifo_reg_2__5_ ( .D(n686), .CLK(clk), .Q(fifo[21]) );
  DFFPOSX1 fifo_reg_2__3_ ( .D(n685), .CLK(clk), .Q(fifo[19]) );
  DFFPOSX1 fifo_reg_2__1_ ( .D(n684), .CLK(clk), .Q(fifo[17]) );
  DFFPOSX1 fifo_reg_2__0_ ( .D(n683), .CLK(clk), .Q(fifo[16]) );
  DFFPOSX1 fifo_reg_2__2_ ( .D(n682), .CLK(clk), .Q(fifo[18]) );
  DFFPOSX1 fifo_reg_2__4_ ( .D(n681), .CLK(clk), .Q(fifo[20]) );
  DFFPOSX1 fifo_reg_2__6_ ( .D(n680), .CLK(clk), .Q(fifo[22]) );
  DFFPOSX1 fifo_reg_1__7_ ( .D(n679), .CLK(clk), .Q(fifo[15]) );
  DFFPOSX1 fifo_reg_1__5_ ( .D(n678), .CLK(clk), .Q(fifo[13]) );
  DFFPOSX1 fifo_reg_1__3_ ( .D(n677), .CLK(clk), .Q(fifo[11]) );
  DFFPOSX1 fifo_reg_1__1_ ( .D(n676), .CLK(clk), .Q(fifo[9]) );
  DFFPOSX1 fifo_reg_1__0_ ( .D(n675), .CLK(clk), .Q(fifo[8]) );
  DFFPOSX1 fifo_reg_1__2_ ( .D(n674), .CLK(clk), .Q(fifo[10]) );
  DFFPOSX1 fifo_reg_1__4_ ( .D(n673), .CLK(clk), .Q(fifo[12]) );
  DFFPOSX1 fifo_reg_1__6_ ( .D(n672), .CLK(clk), .Q(fifo[14]) );
  DFFPOSX1 fifo_reg_0__7_ ( .D(n671), .CLK(clk), .Q(fifo[7]) );
  DFFPOSX1 fifo_reg_0__5_ ( .D(n670), .CLK(clk), .Q(fifo[5]) );
  DFFPOSX1 fifo_reg_0__3_ ( .D(n669), .CLK(clk), .Q(fifo[3]) );
  DFFPOSX1 fifo_reg_0__1_ ( .D(n668), .CLK(clk), .Q(fifo[1]) );
  DFFPOSX1 fifo_reg_0__0_ ( .D(n667), .CLK(clk), .Q(fifo[0]) );
  DFFPOSX1 fifo_reg_0__2_ ( .D(n666), .CLK(clk), .Q(fifo[2]) );
  DFFPOSX1 fifo_reg_0__4_ ( .D(n665), .CLK(clk), .Q(fifo[4]) );
  DFFPOSX1 fifo_reg_0__6_ ( .D(n664), .CLK(clk), .Q(fifo[6]) );
  DFFPOSX1 fifo_reg_7__7_ ( .D(n663), .CLK(clk), .Q(fifo[63]) );
  DFFPOSX1 fifo_reg_7__5_ ( .D(n662), .CLK(clk), .Q(fifo[61]) );
  DFFPOSX1 fifo_reg_7__3_ ( .D(n661), .CLK(clk), .Q(fifo[59]) );
  DFFPOSX1 fifo_reg_7__1_ ( .D(n660), .CLK(clk), .Q(fifo[57]) );
  DFFPOSX1 fifo_reg_7__0_ ( .D(n659), .CLK(clk), .Q(fifo[56]) );
  DFFPOSX1 fifo_reg_7__2_ ( .D(n658), .CLK(clk), .Q(fifo[58]) );
  DFFPOSX1 fifo_reg_7__4_ ( .D(n657), .CLK(clk), .Q(fifo[60]) );
  DFFPOSX1 fifo_reg_7__6_ ( .D(n656), .CLK(clk), .Q(fifo[62]) );
  DFFPOSX1 fifo_reg_6__7_ ( .D(n655), .CLK(clk), .Q(fifo[55]) );
  DFFPOSX1 fifo_reg_6__5_ ( .D(n654), .CLK(clk), .Q(fifo[53]) );
  DFFPOSX1 fifo_reg_6__3_ ( .D(n653), .CLK(clk), .Q(fifo[51]) );
  DFFPOSX1 fifo_reg_6__1_ ( .D(n652), .CLK(clk), .Q(fifo[49]) );
  DFFPOSX1 fifo_reg_6__0_ ( .D(n651), .CLK(clk), .Q(fifo[48]) );
  DFFPOSX1 fifo_reg_6__2_ ( .D(n650), .CLK(clk), .Q(fifo[50]) );
  DFFPOSX1 fifo_reg_6__4_ ( .D(n649), .CLK(clk), .Q(fifo[52]) );
  DFFPOSX1 fifo_reg_6__6_ ( .D(n648), .CLK(clk), .Q(fifo[54]) );
  DFFPOSX1 fifo_reg_5__7_ ( .D(n647), .CLK(clk), .Q(fifo[47]) );
  DFFPOSX1 fifo_reg_5__5_ ( .D(n646), .CLK(clk), .Q(fifo[45]) );
  DFFPOSX1 fifo_reg_5__3_ ( .D(n645), .CLK(clk), .Q(fifo[43]) );
  DFFPOSX1 fifo_reg_5__1_ ( .D(n644), .CLK(clk), .Q(fifo[41]) );
  DFFPOSX1 fifo_reg_5__0_ ( .D(n643), .CLK(clk), .Q(fifo[40]) );
  DFFPOSX1 fifo_reg_5__2_ ( .D(n642), .CLK(clk), .Q(fifo[42]) );
  DFFPOSX1 fifo_reg_5__4_ ( .D(n641), .CLK(clk), .Q(fifo[44]) );
  DFFPOSX1 fifo_reg_5__6_ ( .D(n640), .CLK(clk), .Q(fifo[46]) );
  DFFPOSX1 fifo_reg_4__7_ ( .D(n639), .CLK(clk), .Q(fifo[39]) );
  DFFPOSX1 fifo_reg_4__5_ ( .D(n638), .CLK(clk), .Q(fifo[37]) );
  DFFPOSX1 fifo_reg_4__3_ ( .D(n637), .CLK(clk), .Q(fifo[35]) );
  DFFPOSX1 fifo_reg_4__1_ ( .D(n636), .CLK(clk), .Q(fifo[33]) );
  DFFPOSX1 fifo_reg_4__0_ ( .D(n635), .CLK(clk), .Q(fifo[32]) );
  DFFPOSX1 fifo_reg_4__2_ ( .D(n634), .CLK(clk), .Q(fifo[34]) );
  DFFPOSX1 fifo_reg_4__4_ ( .D(n633), .CLK(clk), .Q(fifo[36]) );
  DFFPOSX1 fifo_reg_4__6_ ( .D(n632), .CLK(clk), .Q(fifo[38]) );
  DFFPOSX1 fifo_reg_15__7_ ( .D(n631), .CLK(clk), .Q(fifo[127]) );
  DFFPOSX1 fifo_reg_15__5_ ( .D(n630), .CLK(clk), .Q(fifo[125]) );
  DFFPOSX1 fifo_reg_15__3_ ( .D(n629), .CLK(clk), .Q(fifo[123]) );
  DFFPOSX1 fifo_reg_15__1_ ( .D(n628), .CLK(clk), .Q(fifo[121]) );
  DFFPOSX1 fifo_reg_15__0_ ( .D(n627), .CLK(clk), .Q(fifo[120]) );
  DFFPOSX1 fifo_reg_15__2_ ( .D(n626), .CLK(clk), .Q(fifo[122]) );
  DFFPOSX1 fifo_reg_15__4_ ( .D(n625), .CLK(clk), .Q(fifo[124]) );
  DFFPOSX1 fifo_reg_15__6_ ( .D(n624), .CLK(clk), .Q(fifo[126]) );
  DFFPOSX1 fifo_reg_14__7_ ( .D(n623), .CLK(clk), .Q(fifo[119]) );
  DFFPOSX1 fifo_reg_14__5_ ( .D(n622), .CLK(clk), .Q(fifo[117]) );
  DFFPOSX1 fifo_reg_14__3_ ( .D(n621), .CLK(clk), .Q(fifo[115]) );
  DFFPOSX1 fifo_reg_14__1_ ( .D(n620), .CLK(clk), .Q(fifo[113]) );
  DFFPOSX1 fifo_reg_14__0_ ( .D(n619), .CLK(clk), .Q(fifo[112]) );
  DFFPOSX1 fifo_reg_14__2_ ( .D(n618), .CLK(clk), .Q(fifo[114]) );
  DFFPOSX1 fifo_reg_14__4_ ( .D(n617), .CLK(clk), .Q(fifo[116]) );
  DFFPOSX1 fifo_reg_14__6_ ( .D(n616), .CLK(clk), .Q(fifo[118]) );
  DFFPOSX1 fifo_reg_13__7_ ( .D(n615), .CLK(clk), .Q(fifo[111]) );
  DFFPOSX1 fifo_reg_13__5_ ( .D(n614), .CLK(clk), .Q(fifo[109]) );
  DFFPOSX1 fifo_reg_13__3_ ( .D(n613), .CLK(clk), .Q(fifo[107]) );
  DFFPOSX1 fifo_reg_13__1_ ( .D(n612), .CLK(clk), .Q(fifo[105]) );
  DFFPOSX1 fifo_reg_13__0_ ( .D(n611), .CLK(clk), .Q(fifo[104]) );
  DFFPOSX1 fifo_reg_13__2_ ( .D(n610), .CLK(clk), .Q(fifo[106]) );
  DFFPOSX1 fifo_reg_13__4_ ( .D(n609), .CLK(clk), .Q(fifo[108]) );
  DFFPOSX1 fifo_reg_13__6_ ( .D(n608), .CLK(clk), .Q(fifo[110]) );
  DFFPOSX1 fifo_reg_12__7_ ( .D(n607), .CLK(clk), .Q(fifo[103]) );
  DFFPOSX1 fifo_reg_12__5_ ( .D(n606), .CLK(clk), .Q(fifo[101]) );
  DFFPOSX1 fifo_reg_12__3_ ( .D(n605), .CLK(clk), .Q(fifo[99]) );
  DFFPOSX1 fifo_reg_12__1_ ( .D(n604), .CLK(clk), .Q(fifo[97]) );
  DFFPOSX1 fifo_reg_12__0_ ( .D(n603), .CLK(clk), .Q(fifo[96]) );
  DFFPOSX1 fifo_reg_12__2_ ( .D(n602), .CLK(clk), .Q(fifo[98]) );
  DFFPOSX1 fifo_reg_12__4_ ( .D(n601), .CLK(clk), .Q(fifo[100]) );
  DFFPOSX1 fifo_reg_12__6_ ( .D(n600), .CLK(clk), .Q(fifo[102]) );
  DFFPOSX1 fifo_reg_11__7_ ( .D(n599), .CLK(clk), .Q(fifo[95]) );
  DFFPOSX1 fifo_reg_11__5_ ( .D(n598), .CLK(clk), .Q(fifo[93]) );
  DFFPOSX1 fifo_reg_11__3_ ( .D(n597), .CLK(clk), .Q(fifo[91]) );
  DFFPOSX1 fifo_reg_11__1_ ( .D(n596), .CLK(clk), .Q(fifo[89]) );
  DFFPOSX1 fifo_reg_11__0_ ( .D(n595), .CLK(clk), .Q(fifo[88]) );
  DFFPOSX1 fifo_reg_11__2_ ( .D(n594), .CLK(clk), .Q(fifo[90]) );
  DFFPOSX1 fifo_reg_11__4_ ( .D(n593), .CLK(clk), .Q(fifo[92]) );
  DFFPOSX1 fifo_reg_11__6_ ( .D(n592), .CLK(clk), .Q(fifo[94]) );
  DFFPOSX1 fifo_reg_10__7_ ( .D(n591), .CLK(clk), .Q(fifo[87]) );
  DFFPOSX1 fifo_reg_10__5_ ( .D(n590), .CLK(clk), .Q(fifo[85]) );
  DFFPOSX1 fifo_reg_10__3_ ( .D(n589), .CLK(clk), .Q(fifo[83]) );
  DFFPOSX1 fifo_reg_10__1_ ( .D(n588), .CLK(clk), .Q(fifo[81]) );
  DFFPOSX1 fifo_reg_10__0_ ( .D(n587), .CLK(clk), .Q(fifo[80]) );
  DFFPOSX1 fifo_reg_10__2_ ( .D(n586), .CLK(clk), .Q(fifo[82]) );
  DFFPOSX1 fifo_reg_10__4_ ( .D(n585), .CLK(clk), .Q(fifo[84]) );
  DFFPOSX1 fifo_reg_10__6_ ( .D(n584), .CLK(clk), .Q(fifo[86]) );
  DFFPOSX1 fifo_reg_9__7_ ( .D(n583), .CLK(clk), .Q(fifo[79]) );
  DFFPOSX1 fifo_reg_9__5_ ( .D(n582), .CLK(clk), .Q(fifo[77]) );
  DFFPOSX1 fifo_reg_9__3_ ( .D(n581), .CLK(clk), .Q(fifo[75]) );
  DFFPOSX1 fifo_reg_9__1_ ( .D(n580), .CLK(clk), .Q(fifo[73]) );
  DFFPOSX1 fifo_reg_9__0_ ( .D(n579), .CLK(clk), .Q(fifo[72]) );
  DFFPOSX1 fifo_reg_9__2_ ( .D(n578), .CLK(clk), .Q(fifo[74]) );
  DFFPOSX1 fifo_reg_9__4_ ( .D(n577), .CLK(clk), .Q(fifo[76]) );
  DFFPOSX1 fifo_reg_9__6_ ( .D(n576), .CLK(clk), .Q(fifo[78]) );
  DFFPOSX1 fifo_reg_8__7_ ( .D(n575), .CLK(clk), .Q(fifo[71]) );
  DFFPOSX1 fifo_reg_8__5_ ( .D(n574), .CLK(clk), .Q(fifo[69]) );
  DFFPOSX1 fifo_reg_8__3_ ( .D(n573), .CLK(clk), .Q(fifo[67]) );
  DFFPOSX1 fifo_reg_8__1_ ( .D(n572), .CLK(clk), .Q(fifo[65]) );
  DFFPOSX1 fifo_reg_8__0_ ( .D(n571), .CLK(clk), .Q(fifo[64]) );
  DFFPOSX1 fifo_reg_8__2_ ( .D(n570), .CLK(clk), .Q(fifo[66]) );
  DFFPOSX1 fifo_reg_8__4_ ( .D(n569), .CLK(clk), .Q(fifo[68]) );
  DFFPOSX1 fifo_reg_8__6_ ( .D(n568), .CLK(clk), .Q(fifo[70]) );
  DFFPOSX1 empty_reg ( .D(n567), .CLK(clk), .Q(empty) );
  DFFPOSX1 full_reg ( .D(n566), .CLK(clk), .Q(full) );
  NAND2X1 U4 ( .A(reset), .B(full), .Y(n365) );
  NAND2X1 U8 ( .A(empty), .B(reset), .Y(n368) );
  FIFO_DW01_inc_0 add_69 ( .A({rd_ptr_4_, n14, n13, n853, n11}), .SUM({n179, 
        n178, n177, n176, n175}) );
  FIFO_DW01_inc_1 add_65 ( .A(wr_ptr), .SUM({n37, n36, n35, n34, n33}) );
  FIFO_DW01_sub_0 sub_38 ( .A(wr_ptr), .B({rd_ptr_4_, n14, n13, n12, n11}), 
        .CI(1'b0), .DIFF(fillcount), .CO(SYNOPSYS_UNCONNECTED_1) );
  INVX2 U355 ( .A(n898), .Y(n906) );
  INVX2 U356 ( .A(n934), .Y(n942) );
  INVX2 U357 ( .A(n945), .Y(n953) );
  AND2X2 U358 ( .A(n731), .B(n727), .Y(n714) );
  AND2X2 U359 ( .A(n734), .B(n731), .Y(n715) );
  AND2X2 U360 ( .A(n916), .B(n733), .Y(n716) );
  AND2X2 U361 ( .A(n731), .B(n733), .Y(n717) );
  AND2X2 U362 ( .A(n916), .B(n732), .Y(n718) );
  AND2X2 U363 ( .A(n731), .B(n732), .Y(n719) );
  AND2X2 U364 ( .A(n734), .B(n916), .Y(n720) );
  AND2X2 U365 ( .A(n734), .B(n987), .Y(n721) );
  AND2X2 U366 ( .A(n734), .B(n996), .Y(n722) );
  AND2X2 U367 ( .A(n732), .B(n987), .Y(n723) );
  AND2X2 U368 ( .A(n732), .B(n996), .Y(n724) );
  AND2X2 U369 ( .A(n733), .B(n987), .Y(n725) );
  AND2X2 U370 ( .A(n733), .B(n996), .Y(n726) );
  AND2X2 U371 ( .A(n1020), .B(wr_ptr[2]), .Y(n727) );
  AND2X2 U372 ( .A(n860), .B(n859), .Y(n728) );
  AND2X2 U373 ( .A(n730), .B(n873), .Y(n731) );
  INVX2 U374 ( .A(n856), .Y(n853) );
  BUFX2 U375 ( .A(n11), .Y(n848) );
  BUFX2 U376 ( .A(n11), .Y(n849) );
  BUFX2 U377 ( .A(n11), .Y(n850) );
  BUFX2 U378 ( .A(n11), .Y(n851) );
  BUFX2 U379 ( .A(n11), .Y(n852) );
  BUFX2 U380 ( .A(n11), .Y(n847) );
  INVX2 U381 ( .A(n175), .Y(n858) );
  INVX2 U382 ( .A(n855), .Y(n854) );
  AND2X1 U383 ( .A(n1037), .B(n1036), .Y(n729) );
  AND2X1 U384 ( .A(n1013), .B(n863), .Y(n730) );
  INVX2 U385 ( .A(n11), .Y(n857) );
  INVX2 U386 ( .A(n12), .Y(n856) );
  INVX2 U387 ( .A(data_in[6]), .Y(n997) );
  INVX2 U388 ( .A(data_in[4]), .Y(n999) );
  INVX2 U389 ( .A(data_in[2]), .Y(n1001) );
  INVX2 U390 ( .A(data_in[0]), .Y(n1003) );
  INVX2 U391 ( .A(data_in[1]), .Y(n1005) );
  INVX2 U392 ( .A(data_in[3]), .Y(n1007) );
  INVX2 U393 ( .A(data_in[5]), .Y(n1009) );
  INVX2 U394 ( .A(data_in[7]), .Y(n1011) );
  INVX2 U395 ( .A(n13), .Y(n855) );
  AND2X1 U396 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .Y(n732) );
  AND2X1 U397 ( .A(wr_ptr[1]), .B(n1018), .Y(n733) );
  NOR2X1 U398 ( .A(wr_ptr[2]), .B(wr_ptr[1]), .Y(n734) );
  MUX2X1 U399 ( .B(n736), .A(n737), .S(n853), .Y(n735) );
  MUX2X1 U400 ( .B(n739), .A(n740), .S(n853), .Y(n738) );
  MUX2X1 U401 ( .B(n742), .A(n743), .S(n853), .Y(n741) );
  MUX2X1 U402 ( .B(n745), .A(n746), .S(n853), .Y(n744) );
  MUX2X1 U403 ( .B(n747), .A(n748), .S(n14), .Y(n174) );
  MUX2X1 U404 ( .B(n750), .A(n751), .S(n853), .Y(n749) );
  MUX2X1 U405 ( .B(n753), .A(n754), .S(n853), .Y(n752) );
  MUX2X1 U406 ( .B(n756), .A(n757), .S(n853), .Y(n755) );
  MUX2X1 U407 ( .B(n759), .A(n760), .S(n853), .Y(n758) );
  MUX2X1 U408 ( .B(n761), .A(n762), .S(n14), .Y(n173) );
  MUX2X1 U409 ( .B(n764), .A(n765), .S(n853), .Y(n763) );
  MUX2X1 U410 ( .B(n767), .A(n768), .S(n853), .Y(n766) );
  MUX2X1 U411 ( .B(n770), .A(n771), .S(n853), .Y(n769) );
  MUX2X1 U412 ( .B(n773), .A(n774), .S(n853), .Y(n772) );
  MUX2X1 U413 ( .B(n775), .A(n776), .S(n14), .Y(n172) );
  MUX2X1 U414 ( .B(n778), .A(n779), .S(n853), .Y(n777) );
  MUX2X1 U415 ( .B(n781), .A(n782), .S(n853), .Y(n780) );
  MUX2X1 U416 ( .B(n784), .A(n785), .S(n853), .Y(n783) );
  MUX2X1 U417 ( .B(n787), .A(n788), .S(n853), .Y(n786) );
  MUX2X1 U418 ( .B(n789), .A(n790), .S(n14), .Y(n171) );
  MUX2X1 U419 ( .B(n792), .A(n793), .S(n853), .Y(n791) );
  MUX2X1 U420 ( .B(n795), .A(n796), .S(n853), .Y(n794) );
  MUX2X1 U421 ( .B(n798), .A(n799), .S(n853), .Y(n797) );
  MUX2X1 U422 ( .B(n801), .A(n802), .S(n853), .Y(n800) );
  MUX2X1 U423 ( .B(n803), .A(n804), .S(n14), .Y(n170) );
  MUX2X1 U424 ( .B(n806), .A(n807), .S(n853), .Y(n805) );
  MUX2X1 U425 ( .B(n809), .A(n810), .S(n853), .Y(n808) );
  MUX2X1 U426 ( .B(n812), .A(n813), .S(n853), .Y(n811) );
  MUX2X1 U427 ( .B(n815), .A(n816), .S(n853), .Y(n814) );
  MUX2X1 U428 ( .B(n817), .A(n818), .S(n14), .Y(n169) );
  MUX2X1 U429 ( .B(n820), .A(n821), .S(n853), .Y(n819) );
  MUX2X1 U430 ( .B(n823), .A(n824), .S(n853), .Y(n822) );
  MUX2X1 U431 ( .B(n826), .A(n827), .S(n853), .Y(n825) );
  MUX2X1 U432 ( .B(n829), .A(n830), .S(n853), .Y(n828) );
  MUX2X1 U433 ( .B(n831), .A(n832), .S(n14), .Y(n168) );
  MUX2X1 U434 ( .B(n834), .A(n835), .S(n853), .Y(n833) );
  MUX2X1 U435 ( .B(n837), .A(n838), .S(n853), .Y(n836) );
  MUX2X1 U436 ( .B(n840), .A(n841), .S(n853), .Y(n839) );
  MUX2X1 U437 ( .B(n843), .A(n844), .S(n853), .Y(n842) );
  MUX2X1 U438 ( .B(n845), .A(n846), .S(n14), .Y(n167) );
  MUX2X1 U439 ( .B(fifo[112]), .A(fifo[120]), .S(n847), .Y(n737) );
  MUX2X1 U440 ( .B(fifo[96]), .A(fifo[104]), .S(n847), .Y(n736) );
  MUX2X1 U441 ( .B(fifo[80]), .A(fifo[88]), .S(n847), .Y(n740) );
  MUX2X1 U442 ( .B(fifo[64]), .A(fifo[72]), .S(n847), .Y(n739) );
  MUX2X1 U443 ( .B(n738), .A(n735), .S(n854), .Y(n748) );
  MUX2X1 U444 ( .B(fifo[48]), .A(fifo[56]), .S(n848), .Y(n743) );
  MUX2X1 U445 ( .B(fifo[32]), .A(fifo[40]), .S(n848), .Y(n742) );
  MUX2X1 U446 ( .B(fifo[16]), .A(fifo[24]), .S(n848), .Y(n746) );
  MUX2X1 U447 ( .B(fifo[0]), .A(fifo[8]), .S(n848), .Y(n745) );
  MUX2X1 U448 ( .B(n744), .A(n741), .S(n854), .Y(n747) );
  MUX2X1 U449 ( .B(fifo[113]), .A(fifo[121]), .S(n848), .Y(n751) );
  MUX2X1 U450 ( .B(fifo[97]), .A(fifo[105]), .S(n848), .Y(n750) );
  MUX2X1 U451 ( .B(fifo[81]), .A(fifo[89]), .S(n848), .Y(n754) );
  MUX2X1 U452 ( .B(fifo[65]), .A(fifo[73]), .S(n848), .Y(n753) );
  MUX2X1 U453 ( .B(n752), .A(n749), .S(n854), .Y(n762) );
  MUX2X1 U454 ( .B(fifo[49]), .A(fifo[57]), .S(n848), .Y(n757) );
  MUX2X1 U455 ( .B(fifo[33]), .A(fifo[41]), .S(n848), .Y(n756) );
  MUX2X1 U456 ( .B(fifo[17]), .A(fifo[25]), .S(n848), .Y(n760) );
  MUX2X1 U457 ( .B(fifo[1]), .A(fifo[9]), .S(n848), .Y(n759) );
  MUX2X1 U458 ( .B(n758), .A(n755), .S(n854), .Y(n761) );
  MUX2X1 U459 ( .B(fifo[114]), .A(fifo[122]), .S(n849), .Y(n765) );
  MUX2X1 U460 ( .B(fifo[98]), .A(fifo[106]), .S(n849), .Y(n764) );
  MUX2X1 U461 ( .B(fifo[82]), .A(fifo[90]), .S(n849), .Y(n768) );
  MUX2X1 U462 ( .B(fifo[66]), .A(fifo[74]), .S(n849), .Y(n767) );
  MUX2X1 U463 ( .B(n766), .A(n763), .S(n854), .Y(n776) );
  MUX2X1 U464 ( .B(fifo[50]), .A(fifo[58]), .S(n849), .Y(n771) );
  MUX2X1 U465 ( .B(fifo[34]), .A(fifo[42]), .S(n849), .Y(n770) );
  MUX2X1 U466 ( .B(fifo[18]), .A(fifo[26]), .S(n849), .Y(n774) );
  MUX2X1 U467 ( .B(fifo[2]), .A(fifo[10]), .S(n849), .Y(n773) );
  MUX2X1 U468 ( .B(n772), .A(n769), .S(n854), .Y(n775) );
  MUX2X1 U469 ( .B(fifo[115]), .A(fifo[123]), .S(n849), .Y(n779) );
  MUX2X1 U470 ( .B(fifo[99]), .A(fifo[107]), .S(n849), .Y(n778) );
  MUX2X1 U471 ( .B(fifo[83]), .A(fifo[91]), .S(n849), .Y(n782) );
  MUX2X1 U472 ( .B(fifo[67]), .A(fifo[75]), .S(n849), .Y(n781) );
  MUX2X1 U473 ( .B(n780), .A(n777), .S(n854), .Y(n790) );
  MUX2X1 U474 ( .B(fifo[51]), .A(fifo[59]), .S(n850), .Y(n785) );
  MUX2X1 U475 ( .B(fifo[35]), .A(fifo[43]), .S(n850), .Y(n784) );
  MUX2X1 U476 ( .B(fifo[19]), .A(fifo[27]), .S(n850), .Y(n788) );
  MUX2X1 U477 ( .B(fifo[3]), .A(fifo[11]), .S(n850), .Y(n787) );
  MUX2X1 U478 ( .B(n786), .A(n783), .S(n854), .Y(n789) );
  MUX2X1 U479 ( .B(fifo[116]), .A(fifo[124]), .S(n850), .Y(n793) );
  MUX2X1 U480 ( .B(fifo[100]), .A(fifo[108]), .S(n850), .Y(n792) );
  MUX2X1 U481 ( .B(fifo[84]), .A(fifo[92]), .S(n850), .Y(n796) );
  MUX2X1 U482 ( .B(fifo[68]), .A(fifo[76]), .S(n850), .Y(n795) );
  MUX2X1 U483 ( .B(n794), .A(n791), .S(n854), .Y(n804) );
  MUX2X1 U484 ( .B(fifo[52]), .A(fifo[60]), .S(n850), .Y(n799) );
  MUX2X1 U485 ( .B(fifo[36]), .A(fifo[44]), .S(n850), .Y(n798) );
  MUX2X1 U486 ( .B(fifo[20]), .A(fifo[28]), .S(n850), .Y(n802) );
  MUX2X1 U487 ( .B(fifo[4]), .A(fifo[12]), .S(n850), .Y(n801) );
  MUX2X1 U488 ( .B(n800), .A(n797), .S(n854), .Y(n803) );
  MUX2X1 U489 ( .B(fifo[117]), .A(fifo[125]), .S(n851), .Y(n807) );
  MUX2X1 U490 ( .B(fifo[101]), .A(fifo[109]), .S(n851), .Y(n806) );
  MUX2X1 U491 ( .B(fifo[85]), .A(fifo[93]), .S(n851), .Y(n810) );
  MUX2X1 U492 ( .B(fifo[69]), .A(fifo[77]), .S(n851), .Y(n809) );
  MUX2X1 U493 ( .B(n808), .A(n805), .S(n854), .Y(n818) );
  MUX2X1 U494 ( .B(fifo[53]), .A(fifo[61]), .S(n851), .Y(n813) );
  MUX2X1 U495 ( .B(fifo[37]), .A(fifo[45]), .S(n851), .Y(n812) );
  MUX2X1 U496 ( .B(fifo[21]), .A(fifo[29]), .S(n851), .Y(n816) );
  MUX2X1 U497 ( .B(fifo[5]), .A(fifo[13]), .S(n851), .Y(n815) );
  MUX2X1 U498 ( .B(n814), .A(n811), .S(n854), .Y(n817) );
  MUX2X1 U499 ( .B(fifo[118]), .A(fifo[126]), .S(n851), .Y(n821) );
  MUX2X1 U500 ( .B(fifo[102]), .A(fifo[110]), .S(n851), .Y(n820) );
  MUX2X1 U501 ( .B(fifo[86]), .A(fifo[94]), .S(n851), .Y(n824) );
  MUX2X1 U502 ( .B(fifo[70]), .A(fifo[78]), .S(n851), .Y(n823) );
  MUX2X1 U503 ( .B(n822), .A(n819), .S(n854), .Y(n832) );
  MUX2X1 U504 ( .B(fifo[54]), .A(fifo[62]), .S(n852), .Y(n827) );
  MUX2X1 U505 ( .B(fifo[38]), .A(fifo[46]), .S(n852), .Y(n826) );
  MUX2X1 U506 ( .B(fifo[22]), .A(fifo[30]), .S(n852), .Y(n830) );
  MUX2X1 U507 ( .B(fifo[6]), .A(fifo[14]), .S(n852), .Y(n829) );
  MUX2X1 U508 ( .B(n828), .A(n825), .S(n854), .Y(n831) );
  MUX2X1 U509 ( .B(fifo[119]), .A(fifo[127]), .S(n852), .Y(n835) );
  MUX2X1 U510 ( .B(fifo[103]), .A(fifo[111]), .S(n852), .Y(n834) );
  MUX2X1 U511 ( .B(fifo[87]), .A(fifo[95]), .S(n852), .Y(n838) );
  MUX2X1 U512 ( .B(fifo[71]), .A(fifo[79]), .S(n852), .Y(n837) );
  MUX2X1 U513 ( .B(n836), .A(n833), .S(n854), .Y(n846) );
  MUX2X1 U514 ( .B(fifo[55]), .A(fifo[63]), .S(n852), .Y(n841) );
  MUX2X1 U515 ( .B(fifo[39]), .A(fifo[47]), .S(n852), .Y(n840) );
  MUX2X1 U516 ( .B(fifo[23]), .A(fifo[31]), .S(n852), .Y(n844) );
  MUX2X1 U517 ( .B(fifo[7]), .A(fifo[15]), .S(n852), .Y(n843) );
  MUX2X1 U518 ( .B(n842), .A(n839), .S(n854), .Y(n845) );
  NOR2X1 U519 ( .A(fillcount[0]), .B(fillcount[1]), .Y(n860) );
  NOR2X1 U520 ( .A(fillcount[2]), .B(fillcount[3]), .Y(n859) );
  NAND2X1 U521 ( .A(fillcount[4]), .B(n728), .Y(n1013) );
  OAI21X1 U522 ( .A(n1013), .B(reset), .C(n365), .Y(n566) );
  INVX2 U523 ( .A(fillcount[4]), .Y(n861) );
  NAND2X1 U524 ( .A(n861), .B(n728), .Y(n1037) );
  OAI21X1 U525 ( .A(n1037), .B(reset), .C(n368), .Y(n567) );
  INVX2 U526 ( .A(fifo[70]), .Y(n865) );
  INVX2 U527 ( .A(put), .Y(n862) );
  NOR2X1 U528 ( .A(reset), .B(n862), .Y(n863) );
  INVX2 U529 ( .A(wr_ptr[0]), .Y(n1022) );
  NAND3X1 U530 ( .A(wr_ptr[3]), .B(n730), .C(n1022), .Y(n864) );
  INVX2 U531 ( .A(n864), .Y(n916) );
  MUX2X1 U532 ( .B(n865), .A(n997), .S(n720), .Y(n568) );
  INVX2 U533 ( .A(fifo[68]), .Y(n866) );
  MUX2X1 U534 ( .B(n866), .A(n999), .S(n720), .Y(n569) );
  INVX2 U535 ( .A(fifo[66]), .Y(n867) );
  MUX2X1 U536 ( .B(n867), .A(n1001), .S(n720), .Y(n570) );
  INVX2 U537 ( .A(fifo[64]), .Y(n868) );
  MUX2X1 U538 ( .B(n868), .A(n1003), .S(n720), .Y(n571) );
  INVX2 U539 ( .A(fifo[65]), .Y(n869) );
  MUX2X1 U540 ( .B(n869), .A(n1005), .S(n720), .Y(n572) );
  INVX2 U541 ( .A(fifo[67]), .Y(n870) );
  MUX2X1 U542 ( .B(n870), .A(n1007), .S(n720), .Y(n573) );
  INVX2 U543 ( .A(fifo[69]), .Y(n871) );
  MUX2X1 U544 ( .B(n871), .A(n1009), .S(n720), .Y(n574) );
  INVX2 U545 ( .A(fifo[71]), .Y(n872) );
  MUX2X1 U546 ( .B(n872), .A(n1011), .S(n720), .Y(n575) );
  INVX2 U547 ( .A(fifo[78]), .Y(n874) );
  AND2X2 U548 ( .A(wr_ptr[0]), .B(wr_ptr[3]), .Y(n873) );
  MUX2X1 U549 ( .B(n874), .A(n997), .S(n715), .Y(n576) );
  INVX2 U550 ( .A(fifo[76]), .Y(n875) );
  MUX2X1 U551 ( .B(n875), .A(n999), .S(n715), .Y(n577) );
  INVX2 U552 ( .A(fifo[74]), .Y(n876) );
  MUX2X1 U553 ( .B(n876), .A(n1001), .S(n715), .Y(n578) );
  INVX2 U554 ( .A(fifo[72]), .Y(n877) );
  MUX2X1 U555 ( .B(n877), .A(n1003), .S(n715), .Y(n579) );
  INVX2 U556 ( .A(fifo[73]), .Y(n878) );
  MUX2X1 U557 ( .B(n878), .A(n1005), .S(n715), .Y(n580) );
  INVX2 U558 ( .A(fifo[75]), .Y(n879) );
  MUX2X1 U559 ( .B(n879), .A(n1007), .S(n715), .Y(n581) );
  INVX2 U560 ( .A(fifo[77]), .Y(n880) );
  MUX2X1 U561 ( .B(n880), .A(n1009), .S(n715), .Y(n582) );
  INVX2 U562 ( .A(fifo[79]), .Y(n881) );
  MUX2X1 U563 ( .B(n881), .A(n1011), .S(n715), .Y(n583) );
  INVX2 U564 ( .A(fifo[86]), .Y(n882) );
  INVX2 U565 ( .A(wr_ptr[2]), .Y(n1018) );
  MUX2X1 U566 ( .B(n882), .A(n997), .S(n716), .Y(n584) );
  INVX2 U567 ( .A(fifo[84]), .Y(n883) );
  MUX2X1 U568 ( .B(n883), .A(n999), .S(n716), .Y(n585) );
  INVX2 U569 ( .A(fifo[82]), .Y(n884) );
  MUX2X1 U570 ( .B(n884), .A(n1001), .S(n716), .Y(n586) );
  INVX2 U571 ( .A(fifo[80]), .Y(n885) );
  MUX2X1 U572 ( .B(n885), .A(n1003), .S(n716), .Y(n587) );
  INVX2 U573 ( .A(fifo[81]), .Y(n886) );
  MUX2X1 U574 ( .B(n886), .A(n1005), .S(n716), .Y(n588) );
  INVX2 U575 ( .A(fifo[83]), .Y(n887) );
  MUX2X1 U576 ( .B(n887), .A(n1007), .S(n716), .Y(n589) );
  INVX2 U577 ( .A(fifo[85]), .Y(n888) );
  MUX2X1 U578 ( .B(n888), .A(n1009), .S(n716), .Y(n590) );
  INVX2 U579 ( .A(fifo[87]), .Y(n889) );
  MUX2X1 U580 ( .B(n889), .A(n1011), .S(n716), .Y(n591) );
  INVX2 U581 ( .A(fifo[94]), .Y(n890) );
  MUX2X1 U582 ( .B(n890), .A(n997), .S(n717), .Y(n592) );
  INVX2 U583 ( .A(fifo[92]), .Y(n891) );
  MUX2X1 U584 ( .B(n891), .A(n999), .S(n717), .Y(n593) );
  INVX2 U585 ( .A(fifo[90]), .Y(n892) );
  MUX2X1 U586 ( .B(n892), .A(n1001), .S(n717), .Y(n594) );
  INVX2 U587 ( .A(fifo[88]), .Y(n893) );
  MUX2X1 U588 ( .B(n893), .A(n1003), .S(n717), .Y(n595) );
  INVX2 U589 ( .A(fifo[89]), .Y(n894) );
  MUX2X1 U590 ( .B(n894), .A(n1005), .S(n717), .Y(n596) );
  INVX2 U591 ( .A(fifo[91]), .Y(n895) );
  MUX2X1 U592 ( .B(n895), .A(n1007), .S(n717), .Y(n597) );
  INVX2 U593 ( .A(fifo[93]), .Y(n896) );
  MUX2X1 U594 ( .B(n896), .A(n1009), .S(n717), .Y(n598) );
  INVX2 U595 ( .A(fifo[95]), .Y(n897) );
  MUX2X1 U596 ( .B(n897), .A(n1011), .S(n717), .Y(n599) );
  INVX2 U597 ( .A(fifo[102]), .Y(n899) );
  INVX2 U598 ( .A(wr_ptr[1]), .Y(n1020) );
  NAND2X1 U599 ( .A(n916), .B(n727), .Y(n898) );
  MUX2X1 U600 ( .B(n899), .A(n997), .S(n906), .Y(n600) );
  INVX2 U601 ( .A(fifo[100]), .Y(n900) );
  MUX2X1 U602 ( .B(n900), .A(n999), .S(n906), .Y(n601) );
  INVX2 U603 ( .A(fifo[98]), .Y(n901) );
  MUX2X1 U604 ( .B(n901), .A(n1001), .S(n906), .Y(n602) );
  INVX2 U605 ( .A(fifo[96]), .Y(n902) );
  MUX2X1 U606 ( .B(n902), .A(n1003), .S(n906), .Y(n603) );
  INVX2 U607 ( .A(fifo[97]), .Y(n903) );
  MUX2X1 U608 ( .B(n903), .A(n1005), .S(n906), .Y(n604) );
  INVX2 U609 ( .A(fifo[99]), .Y(n904) );
  MUX2X1 U610 ( .B(n904), .A(n1007), .S(n906), .Y(n605) );
  INVX2 U611 ( .A(fifo[101]), .Y(n905) );
  MUX2X1 U612 ( .B(n905), .A(n1009), .S(n906), .Y(n606) );
  INVX2 U613 ( .A(fifo[103]), .Y(n907) );
  MUX2X1 U614 ( .B(n907), .A(n1011), .S(n906), .Y(n607) );
  INVX2 U615 ( .A(fifo[110]), .Y(n908) );
  MUX2X1 U616 ( .B(n908), .A(n997), .S(n714), .Y(n608) );
  INVX2 U617 ( .A(fifo[108]), .Y(n909) );
  MUX2X1 U618 ( .B(n909), .A(n999), .S(n714), .Y(n609) );
  INVX2 U619 ( .A(fifo[106]), .Y(n910) );
  MUX2X1 U620 ( .B(n910), .A(n1001), .S(n714), .Y(n610) );
  INVX2 U621 ( .A(fifo[104]), .Y(n911) );
  MUX2X1 U622 ( .B(n911), .A(n1003), .S(n714), .Y(n611) );
  INVX2 U623 ( .A(fifo[105]), .Y(n912) );
  MUX2X1 U624 ( .B(n912), .A(n1005), .S(n714), .Y(n612) );
  INVX2 U625 ( .A(fifo[107]), .Y(n913) );
  MUX2X1 U626 ( .B(n913), .A(n1007), .S(n714), .Y(n613) );
  INVX2 U627 ( .A(fifo[109]), .Y(n914) );
  MUX2X1 U628 ( .B(n914), .A(n1009), .S(n714), .Y(n614) );
  INVX2 U629 ( .A(fifo[111]), .Y(n915) );
  MUX2X1 U630 ( .B(n915), .A(n1011), .S(n714), .Y(n615) );
  INVX2 U631 ( .A(fifo[118]), .Y(n917) );
  MUX2X1 U632 ( .B(n917), .A(n997), .S(n718), .Y(n616) );
  INVX2 U633 ( .A(fifo[116]), .Y(n918) );
  MUX2X1 U634 ( .B(n918), .A(n999), .S(n718), .Y(n617) );
  INVX2 U635 ( .A(fifo[114]), .Y(n919) );
  MUX2X1 U636 ( .B(n919), .A(n1001), .S(n718), .Y(n618) );
  INVX2 U637 ( .A(fifo[112]), .Y(n920) );
  MUX2X1 U638 ( .B(n920), .A(n1003), .S(n718), .Y(n619) );
  INVX2 U639 ( .A(fifo[113]), .Y(n921) );
  MUX2X1 U640 ( .B(n921), .A(n1005), .S(n718), .Y(n620) );
  INVX2 U641 ( .A(fifo[115]), .Y(n922) );
  MUX2X1 U642 ( .B(n922), .A(n1007), .S(n718), .Y(n621) );
  INVX2 U643 ( .A(fifo[117]), .Y(n923) );
  MUX2X1 U644 ( .B(n923), .A(n1009), .S(n718), .Y(n622) );
  INVX2 U645 ( .A(fifo[119]), .Y(n924) );
  MUX2X1 U646 ( .B(n924), .A(n1011), .S(n718), .Y(n623) );
  INVX2 U647 ( .A(fifo[126]), .Y(n925) );
  MUX2X1 U648 ( .B(n925), .A(n997), .S(n719), .Y(n624) );
  INVX2 U649 ( .A(fifo[124]), .Y(n926) );
  MUX2X1 U650 ( .B(n926), .A(n999), .S(n719), .Y(n625) );
  INVX2 U651 ( .A(fifo[122]), .Y(n927) );
  MUX2X1 U652 ( .B(n927), .A(n1001), .S(n719), .Y(n626) );
  INVX2 U653 ( .A(fifo[120]), .Y(n928) );
  MUX2X1 U654 ( .B(n928), .A(n1003), .S(n719), .Y(n627) );
  INVX2 U655 ( .A(fifo[121]), .Y(n929) );
  MUX2X1 U656 ( .B(n929), .A(n1005), .S(n719), .Y(n628) );
  INVX2 U657 ( .A(fifo[123]), .Y(n930) );
  MUX2X1 U658 ( .B(n930), .A(n1007), .S(n719), .Y(n629) );
  INVX2 U659 ( .A(fifo[125]), .Y(n931) );
  MUX2X1 U660 ( .B(n931), .A(n1009), .S(n719), .Y(n630) );
  INVX2 U661 ( .A(fifo[127]), .Y(n932) );
  MUX2X1 U662 ( .B(n932), .A(n1011), .S(n719), .Y(n631) );
  INVX2 U663 ( .A(fifo[38]), .Y(n935) );
  INVX2 U664 ( .A(wr_ptr[3]), .Y(n1025) );
  NAND3X1 U665 ( .A(n1025), .B(n730), .C(n1022), .Y(n933) );
  INVX2 U666 ( .A(n933), .Y(n987) );
  NAND2X1 U667 ( .A(n727), .B(n987), .Y(n934) );
  MUX2X1 U668 ( .B(n935), .A(n997), .S(n942), .Y(n632) );
  INVX2 U669 ( .A(fifo[36]), .Y(n936) );
  MUX2X1 U670 ( .B(n936), .A(n999), .S(n942), .Y(n633) );
  INVX2 U671 ( .A(fifo[34]), .Y(n937) );
  MUX2X1 U672 ( .B(n937), .A(n1001), .S(n942), .Y(n634) );
  INVX2 U673 ( .A(fifo[32]), .Y(n938) );
  MUX2X1 U674 ( .B(n938), .A(n1003), .S(n942), .Y(n635) );
  INVX2 U675 ( .A(fifo[33]), .Y(n939) );
  MUX2X1 U676 ( .B(n939), .A(n1005), .S(n942), .Y(n636) );
  INVX2 U677 ( .A(fifo[35]), .Y(n940) );
  MUX2X1 U678 ( .B(n940), .A(n1007), .S(n942), .Y(n637) );
  INVX2 U679 ( .A(fifo[37]), .Y(n941) );
  MUX2X1 U680 ( .B(n941), .A(n1009), .S(n942), .Y(n638) );
  INVX2 U681 ( .A(fifo[39]), .Y(n943) );
  MUX2X1 U682 ( .B(n943), .A(n1011), .S(n942), .Y(n639) );
  INVX2 U683 ( .A(fifo[46]), .Y(n946) );
  NAND3X1 U684 ( .A(wr_ptr[0]), .B(n730), .C(n1025), .Y(n944) );
  INVX2 U685 ( .A(n944), .Y(n996) );
  NAND2X1 U686 ( .A(n727), .B(n996), .Y(n945) );
  MUX2X1 U687 ( .B(n946), .A(n997), .S(n953), .Y(n640) );
  INVX2 U688 ( .A(fifo[44]), .Y(n947) );
  MUX2X1 U689 ( .B(n947), .A(n999), .S(n953), .Y(n641) );
  INVX2 U690 ( .A(fifo[42]), .Y(n948) );
  MUX2X1 U691 ( .B(n948), .A(n1001), .S(n953), .Y(n642) );
  INVX2 U692 ( .A(fifo[40]), .Y(n949) );
  MUX2X1 U693 ( .B(n949), .A(n1003), .S(n953), .Y(n643) );
  INVX2 U694 ( .A(fifo[41]), .Y(n950) );
  MUX2X1 U695 ( .B(n950), .A(n1005), .S(n953), .Y(n644) );
  INVX2 U696 ( .A(fifo[43]), .Y(n951) );
  MUX2X1 U697 ( .B(n951), .A(n1007), .S(n953), .Y(n645) );
  INVX2 U698 ( .A(fifo[45]), .Y(n952) );
  MUX2X1 U699 ( .B(n952), .A(n1009), .S(n953), .Y(n646) );
  INVX2 U700 ( .A(fifo[47]), .Y(n954) );
  MUX2X1 U701 ( .B(n954), .A(n1011), .S(n953), .Y(n647) );
  INVX2 U702 ( .A(fifo[54]), .Y(n955) );
  MUX2X1 U703 ( .B(n955), .A(n997), .S(n723), .Y(n648) );
  INVX2 U704 ( .A(fifo[52]), .Y(n956) );
  MUX2X1 U705 ( .B(n956), .A(n999), .S(n723), .Y(n649) );
  INVX2 U706 ( .A(fifo[50]), .Y(n957) );
  MUX2X1 U707 ( .B(n957), .A(n1001), .S(n723), .Y(n650) );
  INVX2 U708 ( .A(fifo[48]), .Y(n958) );
  MUX2X1 U709 ( .B(n958), .A(n1003), .S(n723), .Y(n651) );
  INVX2 U710 ( .A(fifo[49]), .Y(n959) );
  MUX2X1 U711 ( .B(n959), .A(n1005), .S(n723), .Y(n652) );
  INVX2 U712 ( .A(fifo[51]), .Y(n960) );
  MUX2X1 U713 ( .B(n960), .A(n1007), .S(n723), .Y(n653) );
  INVX2 U714 ( .A(fifo[53]), .Y(n961) );
  MUX2X1 U715 ( .B(n961), .A(n1009), .S(n723), .Y(n654) );
  INVX2 U716 ( .A(fifo[55]), .Y(n962) );
  MUX2X1 U717 ( .B(n962), .A(n1011), .S(n723), .Y(n655) );
  INVX2 U718 ( .A(fifo[62]), .Y(n963) );
  MUX2X1 U719 ( .B(n963), .A(n997), .S(n724), .Y(n656) );
  INVX2 U720 ( .A(fifo[60]), .Y(n964) );
  MUX2X1 U721 ( .B(n964), .A(n999), .S(n724), .Y(n657) );
  INVX2 U722 ( .A(fifo[58]), .Y(n965) );
  MUX2X1 U723 ( .B(n965), .A(n1001), .S(n724), .Y(n658) );
  INVX2 U724 ( .A(fifo[56]), .Y(n966) );
  MUX2X1 U725 ( .B(n966), .A(n1003), .S(n724), .Y(n659) );
  INVX2 U726 ( .A(fifo[57]), .Y(n967) );
  MUX2X1 U727 ( .B(n967), .A(n1005), .S(n724), .Y(n660) );
  INVX2 U728 ( .A(fifo[59]), .Y(n968) );
  MUX2X1 U729 ( .B(n968), .A(n1007), .S(n724), .Y(n661) );
  INVX2 U730 ( .A(fifo[61]), .Y(n969) );
  MUX2X1 U731 ( .B(n969), .A(n1009), .S(n724), .Y(n662) );
  INVX2 U732 ( .A(fifo[63]), .Y(n970) );
  MUX2X1 U733 ( .B(n970), .A(n1011), .S(n724), .Y(n663) );
  INVX2 U734 ( .A(fifo[6]), .Y(n971) );
  MUX2X1 U735 ( .B(n971), .A(n997), .S(n721), .Y(n664) );
  INVX2 U736 ( .A(fifo[4]), .Y(n972) );
  MUX2X1 U737 ( .B(n972), .A(n999), .S(n721), .Y(n665) );
  INVX2 U738 ( .A(fifo[2]), .Y(n973) );
  MUX2X1 U739 ( .B(n973), .A(n1001), .S(n721), .Y(n666) );
  INVX2 U740 ( .A(fifo[0]), .Y(n974) );
  MUX2X1 U741 ( .B(n974), .A(n1003), .S(n721), .Y(n667) );
  INVX2 U742 ( .A(fifo[1]), .Y(n975) );
  MUX2X1 U743 ( .B(n975), .A(n1005), .S(n721), .Y(n668) );
  INVX2 U744 ( .A(fifo[3]), .Y(n976) );
  MUX2X1 U745 ( .B(n976), .A(n1007), .S(n721), .Y(n669) );
  INVX2 U746 ( .A(fifo[5]), .Y(n977) );
  MUX2X1 U747 ( .B(n977), .A(n1009), .S(n721), .Y(n670) );
  INVX2 U748 ( .A(fifo[7]), .Y(n978) );
  MUX2X1 U749 ( .B(n978), .A(n1011), .S(n721), .Y(n671) );
  INVX2 U750 ( .A(fifo[14]), .Y(n979) );
  MUX2X1 U751 ( .B(n979), .A(n997), .S(n722), .Y(n672) );
  INVX2 U752 ( .A(fifo[12]), .Y(n980) );
  MUX2X1 U753 ( .B(n980), .A(n999), .S(n722), .Y(n673) );
  INVX2 U754 ( .A(fifo[10]), .Y(n981) );
  MUX2X1 U755 ( .B(n981), .A(n1001), .S(n722), .Y(n674) );
  INVX2 U756 ( .A(fifo[8]), .Y(n982) );
  MUX2X1 U757 ( .B(n982), .A(n1003), .S(n722), .Y(n675) );
  INVX2 U758 ( .A(fifo[9]), .Y(n983) );
  MUX2X1 U759 ( .B(n983), .A(n1005), .S(n722), .Y(n676) );
  INVX2 U760 ( .A(fifo[11]), .Y(n984) );
  MUX2X1 U761 ( .B(n984), .A(n1007), .S(n722), .Y(n677) );
  INVX2 U762 ( .A(fifo[13]), .Y(n985) );
  MUX2X1 U763 ( .B(n985), .A(n1009), .S(n722), .Y(n678) );
  INVX2 U764 ( .A(fifo[15]), .Y(n986) );
  MUX2X1 U765 ( .B(n986), .A(n1011), .S(n722), .Y(n679) );
  INVX2 U766 ( .A(fifo[22]), .Y(n988) );
  MUX2X1 U767 ( .B(n988), .A(n997), .S(n725), .Y(n680) );
  INVX2 U768 ( .A(fifo[20]), .Y(n989) );
  MUX2X1 U769 ( .B(n989), .A(n999), .S(n725), .Y(n681) );
  INVX2 U770 ( .A(fifo[18]), .Y(n990) );
  MUX2X1 U771 ( .B(n990), .A(n1001), .S(n725), .Y(n682) );
  INVX2 U772 ( .A(fifo[16]), .Y(n991) );
  MUX2X1 U773 ( .B(n991), .A(n1003), .S(n725), .Y(n683) );
  INVX2 U774 ( .A(fifo[17]), .Y(n992) );
  MUX2X1 U775 ( .B(n992), .A(n1005), .S(n725), .Y(n684) );
  INVX2 U776 ( .A(fifo[19]), .Y(n993) );
  MUX2X1 U777 ( .B(n993), .A(n1007), .S(n725), .Y(n685) );
  INVX2 U778 ( .A(fifo[21]), .Y(n994) );
  MUX2X1 U779 ( .B(n994), .A(n1009), .S(n725), .Y(n686) );
  INVX2 U780 ( .A(fifo[23]), .Y(n995) );
  MUX2X1 U781 ( .B(n995), .A(n1011), .S(n725), .Y(n687) );
  INVX2 U782 ( .A(fifo[30]), .Y(n998) );
  MUX2X1 U783 ( .B(n998), .A(n997), .S(n726), .Y(n688) );
  INVX2 U784 ( .A(fifo[28]), .Y(n1000) );
  MUX2X1 U785 ( .B(n1000), .A(n999), .S(n726), .Y(n689) );
  INVX2 U786 ( .A(fifo[26]), .Y(n1002) );
  MUX2X1 U787 ( .B(n1002), .A(n1001), .S(n726), .Y(n690) );
  INVX2 U788 ( .A(fifo[24]), .Y(n1004) );
  MUX2X1 U789 ( .B(n1004), .A(n1003), .S(n726), .Y(n691) );
  INVX2 U790 ( .A(fifo[25]), .Y(n1006) );
  MUX2X1 U791 ( .B(n1006), .A(n1005), .S(n726), .Y(n692) );
  INVX2 U792 ( .A(fifo[27]), .Y(n1008) );
  MUX2X1 U793 ( .B(n1008), .A(n1007), .S(n726), .Y(n693) );
  INVX2 U794 ( .A(fifo[29]), .Y(n1010) );
  MUX2X1 U795 ( .B(n1010), .A(n1009), .S(n726), .Y(n694) );
  INVX2 U796 ( .A(fifo[31]), .Y(n1012) );
  MUX2X1 U797 ( .B(n1012), .A(n1011), .S(n726), .Y(n695) );
  INVX2 U798 ( .A(reset), .Y(n1028) );
  NAND2X1 U799 ( .A(put), .B(n1013), .Y(n1014) );
  NAND2X1 U800 ( .A(n1028), .B(n1014), .Y(n1026) );
  INVX2 U801 ( .A(wr_ptr[4]), .Y(n1016) );
  NAND2X1 U802 ( .A(n1028), .B(n1026), .Y(n1024) );
  INVX2 U803 ( .A(n37), .Y(n1015) );
  OAI22X1 U804 ( .A(n1026), .B(n1016), .C(n1024), .D(n1015), .Y(n1070) );
  INVX2 U805 ( .A(n35), .Y(n1017) );
  OAI22X1 U806 ( .A(n1026), .B(n1018), .C(n1024), .D(n1017), .Y(n697) );
  INVX2 U807 ( .A(n34), .Y(n1019) );
  OAI22X1 U808 ( .A(n1026), .B(n1020), .C(n1024), .D(n1019), .Y(n698) );
  INVX2 U809 ( .A(n33), .Y(n1021) );
  OAI22X1 U810 ( .A(n1026), .B(n1022), .C(n1024), .D(n1021), .Y(n699) );
  INVX2 U811 ( .A(n36), .Y(n1023) );
  OAI22X1 U812 ( .A(n1026), .B(n1025), .C(n1024), .D(n1023), .Y(n700) );
  NAND2X1 U813 ( .A(get), .B(n1037), .Y(n1027) );
  NAND2X1 U814 ( .A(n1028), .B(n1027), .Y(n1055) );
  INVX2 U815 ( .A(rd_ptr_4_), .Y(n1030) );
  NAND2X1 U816 ( .A(n1028), .B(n1055), .Y(n1054) );
  INVX2 U817 ( .A(n179), .Y(n1029) );
  OAI22X1 U818 ( .A(n1055), .B(n1030), .C(n1054), .D(n1029), .Y(n1069) );
  INVX2 U819 ( .A(n177), .Y(n1031) );
  OAI22X1 U820 ( .A(n1055), .B(n855), .C(n1054), .D(n1031), .Y(n1068) );
  INVX2 U821 ( .A(n176), .Y(n1032) );
  OAI22X1 U822 ( .A(n1055), .B(n856), .C(n1054), .D(n1032), .Y(n1067) );
  INVX2 U823 ( .A(n14), .Y(n1034) );
  INVX2 U824 ( .A(n178), .Y(n1033) );
  OAI22X1 U825 ( .A(n1055), .B(n1034), .C(n1054), .D(n1033), .Y(n1066) );
  INVX2 U826 ( .A(data_out[6]), .Y(n1039) );
  INVX2 U827 ( .A(n168), .Y(n1038) );
  INVX2 U828 ( .A(get), .Y(n1035) );
  NOR2X1 U829 ( .A(reset), .B(n1035), .Y(n1036) );
  MUX2X1 U830 ( .B(n1039), .A(n1038), .S(n729), .Y(n1065) );
  INVX2 U831 ( .A(data_out[4]), .Y(n1041) );
  INVX2 U832 ( .A(n170), .Y(n1040) );
  MUX2X1 U833 ( .B(n1041), .A(n1040), .S(n729), .Y(n1064) );
  INVX2 U834 ( .A(data_out[2]), .Y(n1043) );
  INVX2 U835 ( .A(n172), .Y(n1042) );
  MUX2X1 U836 ( .B(n1043), .A(n1042), .S(n729), .Y(n1063) );
  INVX2 U837 ( .A(data_out[0]), .Y(n1045) );
  INVX2 U838 ( .A(n174), .Y(n1044) );
  MUX2X1 U839 ( .B(n1045), .A(n1044), .S(n729), .Y(n1062) );
  INVX2 U840 ( .A(data_out[1]), .Y(n1047) );
  INVX2 U841 ( .A(n173), .Y(n1046) );
  MUX2X1 U842 ( .B(n1047), .A(n1046), .S(n729), .Y(n1061) );
  INVX2 U843 ( .A(data_out[3]), .Y(n1049) );
  INVX2 U844 ( .A(n171), .Y(n1048) );
  MUX2X1 U845 ( .B(n1049), .A(n1048), .S(n729), .Y(n1060) );
  INVX2 U846 ( .A(data_out[5]), .Y(n1051) );
  INVX2 U847 ( .A(n169), .Y(n1050) );
  MUX2X1 U848 ( .B(n1051), .A(n1050), .S(n729), .Y(n1059) );
  INVX2 U849 ( .A(data_out[7]), .Y(n1053) );
  INVX2 U850 ( .A(n167), .Y(n1052) );
  MUX2X1 U851 ( .B(n1053), .A(n1052), .S(n729), .Y(n1058) );
  OAI22X1 U852 ( .A(n1055), .B(n857), .C(n1054), .D(n858), .Y(n1057) );
endmodule

